magic
tech sky130A
timestamp 1708782296
<< nwell >>
rect -350 -100 1450 400
rect -350 -105 -50 -100
rect 550 -105 850 -100
<< nmos >>
rect -210 -500 -195 -400
rect 90 -500 105 -400
rect 390 -500 405 -400
rect 690 -500 705 -400
rect 990 -500 1005 -400
rect 1290 -500 1305 -400
<< pmos >>
rect -210 -55 -195 145
rect 90 -50 105 150
rect 390 -50 405 150
rect 690 -55 705 145
rect 990 -50 1005 150
rect 1290 -50 1305 150
<< ndiff >>
rect -300 -415 -210 -400
rect -300 -485 -290 -415
rect -225 -485 -210 -415
rect -300 -500 -210 -485
rect -195 -415 -100 -400
rect -195 -485 -180 -415
rect -115 -485 -100 -415
rect -195 -500 -100 -485
rect 0 -415 90 -400
rect 0 -485 15 -415
rect 80 -485 90 -415
rect 0 -500 90 -485
rect 105 -415 200 -400
rect 105 -485 120 -415
rect 185 -485 200 -415
rect 105 -500 200 -485
rect 300 -415 390 -400
rect 300 -485 310 -415
rect 375 -485 390 -415
rect 300 -500 390 -485
rect 405 -415 500 -400
rect 405 -485 420 -415
rect 485 -485 500 -415
rect 405 -500 500 -485
rect 600 -415 690 -400
rect 600 -485 610 -415
rect 675 -485 690 -415
rect 600 -500 690 -485
rect 705 -415 800 -400
rect 705 -485 720 -415
rect 785 -485 800 -415
rect 705 -500 800 -485
rect 900 -415 990 -400
rect 900 -485 915 -415
rect 980 -485 990 -415
rect 900 -500 990 -485
rect 1005 -415 1100 -400
rect 1005 -485 1020 -415
rect 1085 -485 1100 -415
rect 1005 -500 1100 -485
rect 1200 -415 1290 -400
rect 1200 -485 1210 -415
rect 1275 -485 1290 -415
rect 1200 -500 1290 -485
rect 1305 -415 1400 -400
rect 1305 -485 1320 -415
rect 1385 -485 1400 -415
rect 1305 -500 1400 -485
<< pdiff >>
rect -300 130 -225 145
rect -300 -40 -285 130
rect -300 -55 -225 -40
rect -195 140 -100 145
rect -195 130 -120 140
rect -195 -40 -180 130
rect -195 -50 -120 -40
rect -110 -50 -100 140
rect 0 135 75 150
rect 0 -35 15 135
rect 0 -50 75 -35
rect 105 145 200 150
rect 105 135 180 145
rect 105 -35 120 135
rect 105 -45 180 -35
rect 190 -45 200 145
rect 105 -50 200 -45
rect 300 135 375 150
rect 300 -35 315 135
rect 300 -50 375 -35
rect 405 145 500 150
rect 405 135 480 145
rect 405 -35 420 135
rect 405 -45 480 -35
rect 490 -45 500 145
rect 405 -50 500 -45
rect 600 130 675 145
rect 600 -40 615 130
rect -195 -55 -100 -50
rect 600 -55 675 -40
rect 705 140 800 145
rect 705 130 780 140
rect 705 -40 720 130
rect 705 -50 780 -40
rect 790 -50 800 140
rect 900 135 975 150
rect 900 -35 915 135
rect 900 -50 975 -35
rect 1005 145 1100 150
rect 1005 135 1080 145
rect 1005 -35 1020 135
rect 1005 -45 1080 -35
rect 1090 -45 1100 145
rect 1005 -50 1100 -45
rect 1200 135 1275 150
rect 1200 -35 1215 135
rect 1200 -50 1275 -35
rect 1305 145 1400 150
rect 1305 135 1380 145
rect 1305 -35 1320 135
rect 1305 -45 1380 -35
rect 1390 -45 1400 145
rect 1305 -50 1400 -45
rect 705 -55 800 -50
<< ndiffc >>
rect -290 -485 -225 -415
rect -180 -485 -115 -415
rect 15 -485 80 -415
rect 120 -485 185 -415
rect 310 -485 375 -415
rect 420 -485 485 -415
rect 610 -485 675 -415
rect 720 -485 785 -415
rect 915 -485 980 -415
rect 1020 -485 1085 -415
rect 1210 -485 1275 -415
rect 1320 -485 1385 -415
<< pdiffc >>
rect -285 -40 -225 130
rect -180 -40 -120 130
rect 15 -35 75 135
rect 120 -35 180 135
rect 315 -35 375 135
rect 420 -35 480 135
rect 615 -40 675 130
rect 720 -40 780 130
rect 915 -35 975 135
rect 1020 -35 1080 135
rect 1215 -35 1275 135
rect 1320 -35 1380 135
<< psubdiff >>
rect 405 -615 645 -600
rect 405 -730 420 -615
rect 620 -730 645 -615
rect 405 -750 645 -730
<< nsubdiff >>
rect 490 335 690 350
rect 490 280 515 335
rect 655 280 690 335
rect 490 250 690 280
<< psubdiffcont >>
rect 420 -730 620 -615
<< nsubdiffcont >>
rect 515 280 655 335
<< poly >>
rect -210 145 -195 165
rect 90 150 105 170
rect 390 150 405 170
rect 690 145 705 165
rect 990 150 1005 170
rect 1290 150 1305 170
rect -210 -200 -195 -55
rect 90 -200 105 -50
rect 390 -195 405 -50
rect -210 -210 -100 -200
rect -210 -265 -190 -210
rect -105 -265 -100 -210
rect -210 -275 -100 -265
rect -5 -210 105 -200
rect -5 -265 0 -210
rect 85 -265 105 -210
rect -5 -275 105 -265
rect 165 -205 260 -195
rect 165 -260 170 -205
rect 250 -260 260 -205
rect 165 -270 260 -260
rect 295 -205 405 -195
rect 295 -260 305 -205
rect 385 -260 405 -205
rect 525 -175 600 -165
rect 525 -215 535 -175
rect 590 -215 600 -175
rect 525 -225 600 -215
rect 690 -200 705 -55
rect 990 -200 1005 -50
rect 1290 -195 1305 -50
rect 690 -210 800 -200
rect 295 -270 405 -260
rect -210 -400 -195 -275
rect 90 -400 105 -275
rect 390 -400 405 -270
rect 690 -255 710 -210
rect 790 -255 800 -210
rect 690 -265 800 -255
rect 895 -210 1005 -200
rect 895 -255 905 -210
rect 985 -255 1005 -210
rect 895 -265 1005 -255
rect 1065 -205 1160 -195
rect 1065 -250 1070 -205
rect 1150 -250 1160 -205
rect 1065 -260 1160 -250
rect 1195 -205 1305 -195
rect 1195 -250 1205 -205
rect 1285 -250 1305 -205
rect 1195 -260 1305 -250
rect 690 -400 705 -265
rect 990 -400 1005 -265
rect 1290 -400 1305 -260
rect -210 -540 -195 -500
rect 90 -540 105 -500
rect 390 -540 405 -500
rect 690 -540 705 -500
rect 990 -540 1005 -500
rect 1290 -540 1305 -500
<< polycont >>
rect -190 -265 -105 -210
rect 0 -265 85 -210
rect 170 -260 250 -205
rect 305 -260 385 -205
rect 535 -215 590 -175
rect 710 -255 790 -210
rect 905 -255 985 -210
rect 1070 -250 1150 -205
rect 1205 -250 1285 -205
<< pdiffres >>
rect -225 -55 -210 145
rect -120 -50 -110 140
rect 75 -50 90 150
rect 180 -45 190 145
rect 375 -50 390 150
rect 480 -45 490 145
rect 675 -55 690 145
rect 780 -50 790 140
rect 975 -50 990 150
rect 1080 -45 1090 145
rect 1275 -50 1290 150
rect 1380 -45 1390 145
<< locali >>
rect 490 340 690 350
rect -285 335 690 340
rect -285 280 515 335
rect 655 280 965 335
rect -285 140 -230 280
rect 20 145 75 280
rect 490 275 965 280
rect 490 250 690 275
rect 730 225 790 275
rect 620 190 790 225
rect 110 145 175 150
rect -295 130 -215 140
rect -295 -40 -285 130
rect -225 -40 -215 130
rect -295 -50 -215 -40
rect -190 130 -110 140
rect -190 -40 -180 130
rect -115 -40 -110 130
rect -190 -50 -110 -40
rect 5 135 85 145
rect 5 -35 15 135
rect 75 -35 85 135
rect 5 -45 85 -35
rect 110 135 190 145
rect 110 -35 120 135
rect 180 -35 190 135
rect 110 -45 190 -35
rect 305 135 385 145
rect 305 -35 315 135
rect 375 -35 385 135
rect 305 -45 385 -35
rect 410 135 490 145
rect 620 140 680 190
rect 905 145 965 275
rect 410 -35 420 135
rect 480 -35 490 135
rect 410 -45 490 -35
rect 605 130 685 140
rect 605 -40 615 130
rect 675 -40 685 130
rect 115 -195 165 -45
rect 605 -50 685 -40
rect 710 130 790 140
rect 710 -40 720 130
rect 780 -40 790 130
rect 710 -50 790 -40
rect 905 135 985 145
rect 905 -35 915 135
rect 975 -35 985 135
rect 905 -45 985 -35
rect 1010 135 1090 145
rect 1010 -35 1020 135
rect 1080 -35 1090 135
rect 1010 -45 1090 -35
rect 1205 135 1285 145
rect 1205 -35 1215 135
rect 1275 -35 1285 135
rect 1205 -45 1285 -35
rect 1310 135 1390 145
rect 1310 -35 1320 135
rect 1380 -35 1390 135
rect 1310 -45 1390 -35
rect 525 -175 600 -165
rect -195 -210 -100 -200
rect -195 -265 -190 -210
rect -105 -265 -100 -210
rect -195 -275 -100 -265
rect -5 -210 90 -200
rect -5 -265 0 -210
rect 85 -265 90 -210
rect -5 -275 90 -265
rect 115 -205 390 -195
rect 115 -260 170 -205
rect 250 -260 305 -205
rect 385 -260 390 -205
rect 525 -215 535 -175
rect 590 -215 600 -175
rect 1015 -195 1065 -45
rect 525 -225 600 -215
rect 705 -210 800 -200
rect 115 -270 390 -260
rect 705 -255 710 -210
rect 790 -255 800 -210
rect 705 -265 800 -255
rect 895 -210 990 -200
rect 895 -255 905 -210
rect 985 -255 990 -210
rect 895 -265 990 -255
rect 1015 -205 1290 -195
rect 1015 -250 1070 -205
rect 1150 -250 1205 -205
rect 1285 -250 1290 -205
rect 1015 -260 1290 -250
rect 115 -405 165 -270
rect 1015 -405 1065 -260
rect -295 -415 -215 -405
rect -295 -485 -290 -415
rect -225 -485 -215 -415
rect -295 -495 -215 -485
rect -190 -415 -110 -405
rect -190 -485 -180 -415
rect -115 -485 -110 -415
rect -190 -495 -110 -485
rect 10 -415 85 -405
rect 10 -485 15 -415
rect 80 -485 85 -415
rect 10 -495 85 -485
rect 110 -415 190 -405
rect 110 -485 120 -415
rect 185 -485 190 -415
rect 110 -495 190 -485
rect 305 -415 385 -405
rect 305 -485 310 -415
rect 375 -485 385 -415
rect 305 -495 385 -485
rect 410 -415 490 -405
rect 410 -485 420 -415
rect 485 -485 490 -415
rect 410 -495 490 -485
rect 605 -415 685 -405
rect 605 -485 610 -415
rect 675 -485 685 -415
rect 605 -495 685 -485
rect 710 -415 790 -405
rect 710 -485 720 -415
rect 785 -485 790 -415
rect 710 -495 790 -485
rect 910 -415 985 -405
rect 910 -485 915 -415
rect 980 -485 985 -415
rect 910 -495 985 -485
rect 1010 -415 1090 -405
rect 1010 -485 1020 -415
rect 1085 -485 1090 -415
rect 1010 -495 1090 -485
rect 1205 -415 1285 -405
rect 1205 -485 1210 -415
rect 1275 -485 1285 -415
rect 1205 -495 1285 -485
rect 1310 -415 1390 -405
rect 1310 -485 1320 -415
rect 1385 -485 1390 -415
rect 1310 -495 1390 -485
rect 120 -670 185 -495
rect 615 -600 640 -495
rect 405 -615 645 -600
rect 405 -670 420 -615
rect 120 -730 420 -670
rect 620 -670 645 -615
rect 920 -670 980 -495
rect 620 -690 980 -670
rect 1210 -690 1265 -495
rect 620 -730 1265 -690
rect 120 -745 1265 -730
rect 405 -750 645 -745
<< viali >>
rect 515 280 655 335
rect -180 -40 -120 130
rect -120 -40 -115 130
rect 315 -35 375 135
rect 420 -35 480 135
rect 720 -40 780 130
rect 1215 -35 1275 135
rect 1320 -35 1380 135
rect -190 -265 -105 -210
rect 0 -265 85 -210
rect 535 -215 590 -175
rect 710 -255 790 -210
rect 905 -255 985 -210
rect -290 -485 -225 -415
rect -180 -485 -115 -415
rect 310 -485 375 -415
rect 420 -485 485 -415
rect 720 -485 785 -415
rect 1320 -485 1385 -415
<< metal1 >>
rect 490 335 690 350
rect 490 280 515 335
rect 655 280 690 335
rect 490 250 690 280
rect -175 235 440 245
rect -175 225 480 235
rect 1215 225 1275 230
rect -175 195 1275 225
rect -175 140 -115 195
rect 315 145 375 195
rect 440 185 1275 195
rect 440 180 480 185
rect 720 170 1275 185
rect -190 130 -110 140
rect -190 -40 -180 130
rect -115 -40 -110 130
rect -190 -50 -110 -40
rect 305 135 385 145
rect 305 -35 315 135
rect 375 -35 385 135
rect 305 -45 385 -35
rect 410 135 490 145
rect 720 140 765 170
rect 1215 145 1275 170
rect 410 -35 420 135
rect 480 -35 490 135
rect 410 -45 490 -35
rect 710 130 790 140
rect 710 -40 720 130
rect 780 -40 790 130
rect 710 -50 790 -40
rect 1205 135 1285 145
rect 1205 -35 1215 135
rect 1275 -35 1285 135
rect 1205 -45 1285 -35
rect 1310 135 1390 145
rect 1310 -35 1320 135
rect 1380 -35 1390 135
rect 1310 -45 1390 -35
rect 525 -175 600 -165
rect -195 -210 90 -200
rect -195 -265 -190 -210
rect -105 -265 0 -210
rect 85 -265 90 -210
rect 525 -215 535 -175
rect 590 -215 600 -175
rect 525 -225 600 -215
rect 705 -210 990 -200
rect 705 -255 710 -210
rect 790 -255 905 -210
rect 985 -255 990 -210
rect 705 -265 990 -255
rect -195 -275 90 -265
rect -295 -415 -215 -405
rect -295 -485 -290 -415
rect -225 -485 -215 -415
rect -295 -495 -215 -485
rect -190 -415 -110 -405
rect -190 -485 -180 -415
rect -115 -485 -110 -415
rect -190 -495 -110 -485
rect 305 -415 385 -405
rect 305 -485 310 -415
rect 375 -485 385 -415
rect 305 -495 385 -485
rect 410 -415 490 -405
rect 410 -485 420 -415
rect 485 -485 490 -415
rect 410 -495 490 -485
rect 710 -415 790 -405
rect 710 -485 720 -415
rect 785 -485 790 -415
rect 710 -495 790 -485
rect 1310 -415 1390 -405
rect 1310 -485 1320 -415
rect 1385 -485 1390 -415
rect 1310 -495 1390 -485
<< via1 >>
rect 420 -35 480 135
rect 1320 -35 1380 135
rect 535 -215 590 -175
rect -290 -485 -225 -415
rect -180 -485 -115 -415
rect 310 -485 375 -415
rect 420 -485 485 -415
rect 720 -485 785 -415
rect 1320 -485 1385 -415
<< metal2 >>
rect 410 135 490 145
rect 410 -35 420 135
rect 480 -35 490 135
rect 410 -45 490 -35
rect 1310 135 1390 145
rect 1310 -35 1320 135
rect 1380 -35 1390 135
rect 1310 -45 1390 -35
rect 415 -120 485 -45
rect 1320 -120 1390 -45
rect 415 -130 1390 -120
rect -170 -165 1390 -130
rect -170 -170 800 -165
rect -170 -405 -125 -170
rect 430 -405 475 -170
rect 525 -175 600 -170
rect 525 -215 535 -175
rect 590 -215 600 -175
rect 525 -250 600 -215
rect -295 -415 -215 -405
rect -295 -485 -290 -415
rect -225 -485 -215 -415
rect -295 -495 -215 -485
rect -190 -415 -110 -405
rect -190 -485 -180 -415
rect -115 -485 -110 -415
rect -190 -495 -110 -485
rect 305 -415 385 -405
rect 305 -485 310 -415
rect 375 -485 385 -415
rect 305 -495 385 -485
rect 410 -415 490 -405
rect 410 -485 420 -415
rect 485 -485 490 -415
rect 410 -495 490 -485
rect 710 -415 790 -405
rect 710 -485 720 -415
rect 785 -485 790 -415
rect 710 -495 790 -485
rect 1310 -415 1390 -405
rect 1310 -485 1320 -415
rect 1385 -485 1390 -415
rect 1310 -495 1390 -485
<< via2 >>
rect -290 -485 -225 -415
rect 310 -485 375 -415
rect 720 -485 785 -415
rect 1320 -485 1385 -415
<< metal3 >>
rect -285 -360 775 -320
rect -285 -405 -245 -360
rect 730 -405 775 -360
rect -295 -415 -215 -405
rect -295 -485 -290 -415
rect -225 -485 -215 -415
rect -295 -495 -215 -485
rect 305 -415 385 -405
rect 305 -485 310 -415
rect 375 -485 385 -415
rect 305 -495 385 -485
rect 710 -415 790 -405
rect 710 -485 720 -415
rect 785 -485 790 -415
rect 710 -495 790 -485
rect 1310 -415 1390 -405
rect 1310 -485 1320 -415
rect 1385 -485 1390 -415
rect 1310 -495 1390 -485
rect 315 -570 375 -495
rect 1330 -570 1385 -495
rect 315 -630 1385 -570
<< labels >>
rlabel metal2 570 -240 570 -240 1 c
port 1 n
rlabel metal1 -50 -240 -50 -240 1 a
port 2 n
rlabel metal1 840 -235 840 -235 1 b
port 3 n
rlabel locali 715 -715 715 -715 1 gnd
port 4 n
rlabel locali 470 310 470 310 1 vdd
port 5 n
<< end >>
