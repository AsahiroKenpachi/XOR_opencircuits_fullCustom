* SPICE3 file created from new4.ext - technology: sky130A


X0 a_300_n500# a_1005_n500# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.95 pd=3.9 as=0.9 ps=3.8 w=1 l=0.15
X1 c a_105_n500# a_n195_n55# vdd sky130_fd_pr__pfet_01v8 ad=1.3 pd=5.3 as=1.3 ps=5.3 w=2 l=0.15
X2 a_n195_n55# b vdd vdd sky130_fd_pr__pfet_01v8 ad=1.3 pd=5.3 as=1.3 ps=5.3 w=2 l=0.15
X3 c a_105_n500# a_300_n500# gnd sky130_fd_pr__nfet_01v8 ad=0.95 pd=3.9 as=0.9 ps=3.8 w=1 l=0.15
X4 a_1005_n500# b vdd vdd sky130_fd_pr__pfet_01v8 ad=1.3 pd=5.3 as=1.3 ps=5.3 w=2 l=0.15
X5 a_105_n500# a vdd vdd sky130_fd_pr__pfet_01v8 ad=1.3 pd=5.3 as=1.3 ps=5.3 w=2 l=0.15
X6 a_n195_n55# a vdd vdd sky130_fd_pr__pfet_01v8 ad=1.3 pd=5.3 as=1.3 ps=5.3 w=2 l=0.15
X7 c a_1005_n500# a_n195_n55# vdd sky130_fd_pr__pfet_01v8 ad=1.3 pd=5.3 as=1.3 ps=5.3 w=2 l=0.15
X8 a_n300_n500# b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.95 pd=3.9 as=0.9 ps=3.8 w=1 l=0.15
X9 a_105_n500# a gnd gnd sky130_fd_pr__nfet_01v8 ad=0.95 pd=3.9 as=0.9 ps=3.8 w=1 l=0.15
X10 c a a_n300_n500# gnd sky130_fd_pr__nfet_01v8 ad=0.95 pd=3.9 as=0.9 ps=3.8 w=1 l=0.15
X11 a_1005_n500# b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.95 pd=3.9 as=0.9 ps=3.8 w=1 l=0.15


